module display_controller(num, num_on_display);

input logic[9:0] num;
output logic[20:0] num_on_display;

logic[3:0] num0 = 0;
logic[3:0] num1 = 0;
logic[3:0] num2 = 0;

endmodule
